module F1VU9PWrapper(
  input          clk_main_a0,
  input          tck,
  input          tms,
  input          tdi,
  output         tdo,
  input  [15:0]  sh_cl_status_vdip,
  output [15:0]  cl_sh_status_vled,
  inout  [17:0]  M_D_DQS_DN,
  inout  [17:0]  M_D_DQS_DP,
  inout  [7:0]   M_D_ECC,
  inout  [63:0]  M_D_DQ,
  inout  [17:0]  M_B_DQS_DN,
  inout  [17:0]  M_B_DQS_DP,
  inout  [7:0]   M_B_ECC,
  inout  [63:0]  M_B_DQ,
  inout  [17:0]  M_A_DQS_DN,
  inout  [17:0]  M_A_DQS_DP,
  inout  [7:0]   M_A_ECC,
  inout  [63:0]  M_A_DQ,
  output [7:0]   ddr_sh_stat_int2,
  output [31:0]  ddr_sh_stat_rdata2,
  output         ddr_sh_stat_ack2,
  input  [31:0]  sh_ddr_stat_wdata2,
  input          sh_ddr_stat_rd2,
  input          sh_ddr_stat_wr2,
  input  [7:0]   sh_ddr_stat_addr2,
  output [7:0]   ddr_sh_stat_int1,
  output [31:0]  ddr_sh_stat_rdata1,
  output         ddr_sh_stat_ack1,
  input  [31:0]  sh_ddr_stat_wdata1,
  input          sh_ddr_stat_rd1,
  input          sh_ddr_stat_wr1,
  input  [7:0]   sh_ddr_stat_addr1,
  output [7:0]   ddr_sh_stat_int0,
  output [31:0]  ddr_sh_stat_rdata0,
  output         ddr_sh_stat_ack0,
  input  [31:0]  sh_ddr_stat_wdata0,
  input          sh_ddr_stat_rd0,
  input          sh_ddr_stat_wr0,
  input  [7:0]   sh_ddr_stat_addr0,
  output         cl_RST_DIMM_D_N,
  output         M_D_PAR,
  output [0:0]   M_D_CLK_DP,
  output [0:0]   M_D_CLK_DN,
  output [0:0]   M_D_CS_N,
  output [0:0]   M_D_ODT,
  output [0:0]   M_D_CKE,
  output [1:0]   M_D_BG,
  output [1:0]   M_D_BA,
  output [16:0]  M_D_MA,
  output         M_D_ACT_N,
  input          CLK_300M_DIMM3_DN,
  input          CLK_300M_DIMM3_DP,
  output         cl_RST_DIMM_B_N,
  output         M_B_PAR,
  output [0:0]   M_B_CLK_DP,
  output [0:0]   M_B_CLK_DN,
  output [0:0]   M_B_CS_N,
  output [0:0]   M_B_ODT,
  output [0:0]   M_B_CKE,
  output [1:0]   M_B_BG,
  output [1:0]   M_B_BA,
  output [16:0]  M_B_MA,
  output         M_B_ACT_N,
  input          CLK_300M_DIMM1_DN,
  input          CLK_300M_DIMM1_DP,
  output         cl_RST_DIMM_A_N,
  output         M_A_PAR,
  output [0:0]   M_A_CLK_DP,
  output [0:0]   M_A_CLK_DN,
  output [0:0]   M_A_CS_N,
  output [0:0]   M_A_ODT,
  output [0:0]   M_A_CKE,
  output [1:0]   M_A_BG,
  output [1:0]   M_A_BA,
  output [16:0]  M_A_MA,
  output         M_A_ACT_N,
  input          CLK_300M_DIMM0_DN,
  input          CLK_300M_DIMM0_DP,
  input          rst_main_n,
  output [31:0]  cl_sh_id0,
  output [31:0]  cl_sh_id1,
  input          clk_extra_a1,
  input          clk_extra_a2,
  input          clk_extra_a3,
  input          clk_extra_b0,
  input          clk_extra_b1,
  input          clk_extra_c0,
  input          clk_extra_c1,
  input          kernel_rst_n,
  input          sh_cl_flr_assert,
  output         cl_sh_flr_done,
  output [31:0]  cl_sh_status0,
  output [31:0]  cl_sh_status1,
  input  [31:0]  sh_cl_ctl0,
  input  [31:0]  sh_cl_ctl1,
  input  [1:0]   sh_cl_pwr_state,
  output         cl_sh_dma_wr_full,
  output         cl_sh_dma_rd_full,
  output [15:0]  cl_sh_pcim_awid,
  output [63:0]  cl_sh_pcim_awaddr,
  output [7:0]   cl_sh_pcim_awlen,
  output [2:0]   cl_sh_pcim_awsize,
  output [18:0]  cl_sh_pcim_awuser,
  output         cl_sh_pcim_awvalid,
  input          sh_cl_pcim_awready,
  output [511:0] cl_sh_pcim_wdata,
  output [63:0]  cl_sh_pcim_wstrb,
  output         cl_sh_pcim_wlast,
  output         cl_sh_pcim_wvalid,
  input          sh_cl_pcim_wready,
  input  [15:0]  sh_cl_pcim_bid,
  input  [1:0]   sh_cl_pcim_bresp,
  input          sh_cl_pcim_bvalid,
  output         cl_sh_pcim_bready,
  output [15:0]  cl_sh_pcim_arid,
  output [63:0]  cl_sh_pcim_araddr,
  output [7:0]   cl_sh_pcim_arlen,
  output [2:0]   cl_sh_pcim_arsize,
  output [18:0]  cl_sh_pcim_aruser,
  output         cl_sh_pcim_arvalid,
  input          sh_cl_pcim_arready,
  input  [15:0]  sh_cl_pcim_rid,
  input  [511:0] sh_cl_pcim_rdata,
  input  [1:0]   sh_cl_pcim_rresp,
  input          sh_cl_pcim_rlast,
  input          sh_cl_pcim_rvalid,
  output         cl_sh_pcim_rready,
  input  [1:0]   cfg_max_payload,
  input  [2:0]   cfg_max_read_req,
  output [15:0]  cl_sh_ddr_awid,
  output [63:0]  cl_sh_ddr_awaddr,
  output [7:0]   cl_sh_ddr_awlen,
  output [2:0]   cl_sh_ddr_awsize,
  output [1:0]   cl_sh_ddr_awburst,
  output         cl_sh_ddr_awvalid,
  input          sh_cl_ddr_awready,
  output [15:0]  cl_sh_ddr_wid,
  output [511:0] cl_sh_ddr_wdata,
  output [63:0]  cl_sh_ddr_wstrb,
  output         cl_sh_ddr_wlast,
  output         cl_sh_ddr_wvalid,
  input          sh_cl_ddr_wready,
  input  [15:0]  sh_cl_ddr_bid,
  input  [1:0]   sh_cl_ddr_bresp,
  input          sh_cl_ddr_bvalid,
  output         cl_sh_ddr_bready,
  output [15:0]  cl_sh_ddr_arid,
  output [63:0]  cl_sh_ddr_araddr,
  output [7:0]   cl_sh_ddr_arlen,
  output [2:0]   cl_sh_ddr_arsize,
  output [1:0]   cl_sh_ddr_arburst,
  output         cl_sh_ddr_arvalid,
  input          sh_cl_ddr_arready,
  input  [15:0]  sh_cl_ddr_rid,
  input  [511:0] sh_cl_ddr_rdata,
  input  [1:0]   sh_cl_ddr_rresp,
  input          sh_cl_ddr_rlast,
  input          sh_cl_ddr_rvalid,
  output         cl_sh_ddr_rready,
  input          sh_cl_ddr_is_ready,
  output [15:0]  cl_sh_apppf_irq_req,
  input  [15:0]  sh_cl_apppf_irq_ack,
  input  [5:0]   sh_cl_dma_pcis_awid,
  input  [63:0]  sh_cl_dma_pcis_awaddr,
  input  [7:0]   sh_cl_dma_pcis_awlen,
  input  [2:0]   sh_cl_dma_pcis_awsize,
  input          sh_cl_dma_pcis_awvalid,
  output         cl_sh_dma_pcis_awready,
  input  [511:0] sh_cl_dma_pcis_wdata,
  input  [63:0]  sh_cl_dma_pcis_wstrb,
  input          sh_cl_dma_pcis_wlast,
  input          sh_cl_dma_pcis_wvalid,
  output         cl_sh_dma_pcis_wready,
  output [5:0]   cl_sh_dma_pcis_bid,
  output [1:0]   cl_sh_dma_pcis_bresp,
  output         cl_sh_dma_pcis_bvalid,
  input          sh_cl_dma_pcis_bready,
  input  [5:0]   sh_cl_dma_pcis_arid,
  input  [63:0]  sh_cl_dma_pcis_araddr,
  input  [7:0]   sh_cl_dma_pcis_arlen,
  input  [2:0]   sh_cl_dma_pcis_arsize,
  input          sh_cl_dma_pcis_arvalid,
  output         cl_sh_dma_pcis_arready,
  output [5:0]   cl_sh_dma_pcis_rid,
  output [511:0] cl_sh_dma_pcis_rdata,
  output [1:0]   cl_sh_dma_pcis_rresp,
  output         cl_sh_dma_pcis_rlast,
  output         cl_sh_dma_pcis_rvalid,
  input          sh_cl_dma_pcis_rready,
  input          sda_cl_awvalid,
  input  [31:0]  sda_cl_awaddr,
  output         cl_sda_awready,
  input          sda_cl_wvalid,
  input  [31:0]  sda_cl_wdata,
  input  [3:0]   sda_cl_wstrb,
  output         cl_sda_wready,
  output         cl_sda_bvalid,
  output [1:0]   cl_sda_bresp,
  input          sda_cl_bready,
  input          sda_cl_arvalid,
  input  [31:0]  sda_cl_araddr,
  output         cl_sda_arready,
  output         cl_sda_rvalid,
  output [31:0]  cl_sda_rdata,
  output [1:0]   cl_sda_rresp,
  input          sda_cl_rready,
  input          sh_ocl_awvalid,
  input  [31:0]  sh_ocl_awaddr,
  output         ocl_sh_awready,
  input          sh_ocl_wvalid,
  input  [31:0]  sh_ocl_wdata,
  input  [3:0]   sh_ocl_wstrb,
  output         ocl_sh_wready,
  output         ocl_sh_bvalid,
  output [1:0]   ocl_sh_bresp,
  input          sh_ocl_bready,
  input          sh_ocl_arvalid,
  input  [31:0]  sh_ocl_araddr,
  output         ocl_sh_arready,
  output         ocl_sh_rvalid,
  output [31:0]  ocl_sh_rdata,
  output [1:0]   ocl_sh_rresp,
  input          sh_ocl_rready,
  input          sh_bar1_awvalid,
  input  [31:0]  sh_bar1_awaddr,
  output         bar1_sh_awready,
  input          sh_bar1_wvalid,
  input  [31:0]  sh_bar1_wdata,
  input  [3:0]   sh_bar1_wstrb,
  output         bar1_sh_wready,
  output         bar1_sh_bvalid,
  output [1:0]   bar1_sh_bresp,
  input          sh_bar1_bready,
  input          sh_bar1_arvalid,
  input  [31:0]  sh_bar1_araddr,
  output         bar1_sh_arready,
  output         bar1_sh_rvalid,
  output [31:0]  bar1_sh_rdata,
  output [1:0]   bar1_sh_rresp,
  input          sh_bar1_rready,
  input          drck,
  input          shift,
  input          update,
  input          sel,
  input          runtest,
  input          reset,
  input          capture,
  input          bscanid_en,
  input  [63:0]  sh_cl_glcount0,
  input  [63:0]  sh_cl_glcount1
);
	wire M_A_CKE0;
	wire M_A_ODT0;
	wire M_A_CS_N0;
	wire M_A_CLK_DN0;
	wire M_A_CLK_DP0;
	wire M_B_CKE0;
	wire M_B_ODT0;
	wire M_B_CS_N0;
	wire M_B_CLK_DN0;
	wire M_B_CLK_DP0;
	wire M_D_CKE0;
	wire M_D_ODT0;
	wire M_D_CS_N0;
	wire M_D_CLK_DN0;
	wire M_D_CLK_DP0;
	assign M_A_CKE[0] = M_A_CKE0;
	assign M_A_ODT[0] = M_A_ODT0;
	assign M_A_CS_N[0] = M_A_CS_N0;
	assign M_A_CLK_DN[0] = M_A_CKE0;
	assign M_A_CLK_DP[0] = M_A_CKE0;
	assign M_B_CKE[0] = M_B_CKE0;
	assign M_B_ODT[0] = M_B_ODT0;
	assign M_B_CS_N[0] = M_B_CS_N0;
	assign M_B_CLK_DN[0] = M_B_CKE0;
	assign M_B_CLK_DP[0] = M_B_CKE0;
	assign M_D_CKE[0] = M_D_CKE0;
	assign M_D_ODT[0] = M_D_ODT0;
	assign M_D_CS_N[0] = M_D_CS_N0;
	assign M_D_CLK_DN[0] = M_D_CKE0;
	assign M_D_CLK_DP[0] = M_D_CKE0;
	F1VU9PShell shell (
	  .clk_main_a0(clk_main_a0),
    .tck(tck),
    .tms(tms),
    .tdi(tdi),
    .tdo(tdo),
    .sh_cl_status_vdip(sh_cl_status_vdip),
    .cl_sh_status_vled(cl_sh_status_vled),
    .M_D_DQS_DN(M_D_DQS_DN),
    .M_D_DQS_DP(M_D_DQS_DP),
    .M_D_ECC(M_D_ECC),
    .M_D_DQ(M_D_DQ),
    .M_B_DQS_DN(M_B_DQS_DN),
    .M_B_DQS_DP(M_B_DQS_DP),
    .M_B_ECC(M_B_ECC),
    .M_B_DQ(M_B_DQ),
    .M_A_DQS_DN(M_A_DQS_DN),
    .M_A_DQS_DP(M_A_DQS_DP),
    .M_A_ECC(M_A_ECC),
    .M_A_DQ(M_A_DQ),
    .ddr_sh_stat_int2(ddr_sh_stat_int2),
    .ddr_sh_stat_rdata2(ddr_sh_stat_rdata2),
    .ddr_sh_stat_ack2(ddr_sh_stat_ack2),
    .sh_ddr_stat_wdata2(sh_ddr_stat_wdata2),
    .sh_ddr_stat_rd2(sh_ddr_stat_rd2),
    .sh_ddr_stat_wr2(sh_ddr_stat_wr2),
    .sh_ddr_stat_addr2(sh_ddr_stat_addr2),
    .ddr_sh_stat_int1(ddr_sh_stat_int1),
    .ddr_sh_stat_rdata1(ddr_sh_stat_rdata1),
    .ddr_sh_stat_ack1(ddr_sh_stat_ack1),
    .sh_ddr_stat_wdata1(sh_ddr_stat_wdata1),
    .sh_ddr_stat_rd1(sh_ddr_stat_rd1),
    .sh_ddr_stat_wr1(sh_ddr_stat_wr1),
    .sh_ddr_stat_addr1(sh_ddr_stat_addr1),
    .ddr_sh_stat_int0(ddr_sh_stat_int0),
    .ddr_sh_stat_rdata0(ddr_sh_stat_rdata0),
    .ddr_sh_stat_ack0(ddr_sh_stat_ack0),
    .sh_ddr_stat_wdata0(sh_ddr_stat_wdata0),
    .sh_ddr_stat_rd0(sh_ddr_stat_rd0),
    .sh_ddr_stat_wr0(sh_ddr_stat_wr0),
    .sh_ddr_stat_addr0(sh_ddr_stat_addr0),
    .cl_RST_DIMM_D_N(cl_RST_DIMM_D_N),
    .M_D_PAR(M_D_PAR),
    .M_D_CLK_DP(M_D_CLK_DP0),
    .M_D_CLK_DN(M_D_CLK_DN0),
    .M_D_CS_N(M_D_CS_N0),
    .M_D_ODT(M_D_ODT0),
    .M_D_CKE(M_D_CKE0),
    .M_D_BG(M_D_BG),
    .M_D_BA(M_D_BA),
    .M_D_MA(M_D_MA),
    .M_D_ACT_N(M_D_ACT_N),
    .CLK_300M_DIMM3_DN(CLK_300M_DIMM3_DN),
    .CLK_300M_DIMM3_DP(CLK_300M_DIMM3_DP),
    .cl_RST_DIMM_B_N(cl_RST_DIMM_B_N),
    .M_B_PAR(M_B_PAR),
    .M_B_CLK_DP(M_B_CLK_DP0),
    .M_B_CLK_DN(M_B_CLK_DN0),
    .M_B_CS_N(M_B_CS_N0),
    .M_B_ODT(M_B_ODT0),
    .M_B_CKE(M_B_CKE0),
    .M_B_BG(M_B_BG),
    .M_B_BA(M_B_BA),
    .M_B_MA(M_B_MA),
    .M_B_ACT_N(M_B_ACT_N),
    .CLK_300M_DIMM1_DN(CLK_300M_DIMM1_DN),
    .CLK_300M_DIMM1_DP(CLK_300M_DIMM1_DP),
    .cl_RST_DIMM_A_N(cl_RST_DIMM_A_N),
    .M_A_PAR(M_A_PAR),
    .M_A_CLK_DP(M_A_CLK_DP0),
    .M_A_CLK_DN(M_A_CLK_DN0),
    .M_A_CS_N(M_A_CS_N0),
    .M_A_ODT(M_A_ODT0),
    .M_A_CKE(M_A_CKE0),
    .M_A_BG(M_A_BG),
    .M_A_BA(M_A_BA),
    .M_A_MA(M_A_MA),
    .M_A_ACT_N(M_A_ACT_N),
    .CLK_300M_DIMM0_DN(CLK_300M_DIMM0_DN),
    .CLK_300M_DIMM0_DP(CLK_300M_DIMM0_DP),
    .rst_main_n(rst_main_n),
    .cl_sh_id0(cl_sh_id0),
    .cl_sh_id1(cl_sh_id1),
    .clk_extra_a1(clk_extra_a1),
    .clk_extra_a2(clk_extra_a2),
    .clk_extra_a3(clk_extra_a3),
    .clk_extra_b0(clk_extra_b0),
    .clk_extra_b1(clk_extra_b1),
    .clk_extra_c0(clk_extra_c0),
    .clk_extra_c1(clk_extra_c1),
    .kernel_rst_n(kernel_rst_n),
    .sh_cl_flr_assert(sh_cl_flr_assert),
    .cl_sh_flr_done(cl_sh_flr_done),
    .cl_sh_status0(cl_sh_status0),
    .cl_sh_status1(cl_sh_status1),
    .sh_cl_ctl0(sh_cl_ctl0),
    .sh_cl_ctl1(sh_cl_ctl1),
    .sh_cl_pwr_state(sh_cl_pwr_state),
    .cl_sh_dma_wr_full(cl_sh_dma_wr_full),
    .cl_sh_dma_rd_full(cl_sh_dma_rd_full),
    .cl_sh_pcim_awid(cl_sh_pcim_awid),
    .cl_sh_pcim_awaddr(cl_sh_pcim_awaddr),
    .cl_sh_pcim_awlen(cl_sh_pcim_awlen),
    .cl_sh_pcim_awsize(cl_sh_pcim_awsize),
    .cl_sh_pcim_awuser(cl_sh_pcim_awuser),
    .cl_sh_pcim_awvalid(cl_sh_pcim_awvalid),
    .sh_cl_pcim_awready(sh_cl_pcim_awready),
    .cl_sh_pcim_wdata(cl_sh_pcim_wdata),
    .cl_sh_pcim_wstrb(cl_sh_pcim_wstrb),
    .cl_sh_pcim_wlast(cl_sh_pcim_wlast),
    .cl_sh_pcim_wvalid(cl_sh_pcim_wvalid),
    .sh_cl_pcim_wready(sh_cl_pcim_wready),
    .sh_cl_pcim_bid(sh_cl_pcim_bid),
    .sh_cl_pcim_bresp(sh_cl_pcim_bresp),
    .sh_cl_pcim_bvalid(sh_cl_pcim_bvalid),
    .cl_sh_pcim_bready(cl_sh_pcim_bready),
    .cl_sh_pcim_arid(cl_sh_pcim_arid),
    .cl_sh_pcim_araddr(cl_sh_pcim_araddr),
    .cl_sh_pcim_arlen(cl_sh_pcim_arlen),
    .cl_sh_pcim_arsize(cl_sh_pcim_arsize),
    .cl_sh_pcim_aruser(cl_sh_pcim_aruser),
    .cl_sh_pcim_arvalid(cl_sh_pcim_arvalid),
    .sh_cl_pcim_arready(sh_cl_pcim_arready),
    .sh_cl_pcim_rid(sh_cl_pcim_rid),
    .sh_cl_pcim_rdata(sh_cl_pcim_rdata),
    .sh_cl_pcim_rresp(sh_cl_pcim_rresp),
    .sh_cl_pcim_rlast(sh_cl_pcim_rlast),
    .sh_cl_pcim_rvalid(sh_cl_pcim_rvalid),
    .cl_sh_pcim_rready(cl_sh_pcim_rready),
    .cfg_max_payload(cfg_max_payload),
    .cfg_max_read_req(cfg_max_read_req),
    .cl_sh_ddr_awid(cl_sh_ddr_awid),
    .cl_sh_ddr_awaddr(cl_sh_ddr_awaddr),
    .cl_sh_ddr_awlen(cl_sh_ddr_awlen),
    .cl_sh_ddr_awsize(cl_sh_ddr_awsize),
    .cl_sh_ddr_awburst(cl_sh_ddr_awburst),
    .cl_sh_ddr_awvalid(cl_sh_ddr_awvalid),
    .sh_cl_ddr_awready(sh_cl_ddr_awready),
    .cl_sh_ddr_wid(cl_sh_ddr_wid),
    .cl_sh_ddr_wdata(cl_sh_ddr_wdata),
    .cl_sh_ddr_wstrb(cl_sh_ddr_wstrb),
    .cl_sh_ddr_wlast(cl_sh_ddr_wlast),
    .cl_sh_ddr_wvalid(cl_sh_ddr_wvalid),
    .sh_cl_ddr_wready(sh_cl_ddr_wready),
    .sh_cl_ddr_bid(sh_cl_ddr_bid),
    .sh_cl_ddr_bresp(sh_cl_ddr_bresp),
    .sh_cl_ddr_bvalid(sh_cl_ddr_bvalid),
    .cl_sh_ddr_bready(cl_sh_ddr_bready),
    .cl_sh_ddr_arid(cl_sh_ddr_arid),
    .cl_sh_ddr_araddr(cl_sh_ddr_araddr),
    .cl_sh_ddr_arlen(cl_sh_ddr_arlen),
    .cl_sh_ddr_arsize(cl_sh_ddr_arsize),
    .cl_sh_ddr_arburst(cl_sh_ddr_arburst),
    .cl_sh_ddr_arvalid(cl_sh_ddr_arvalid),
    .sh_cl_ddr_arready(sh_cl_ddr_arready),
    .sh_cl_ddr_rid(sh_cl_ddr_rid),
    .sh_cl_ddr_rdata(sh_cl_ddr_rdata),
    .sh_cl_ddr_rresp(sh_cl_ddr_rresp),
    .sh_cl_ddr_rlast(sh_cl_ddr_rlast),
    .sh_cl_ddr_rvalid(sh_cl_ddr_rvalid),
    .cl_sh_ddr_rready(cl_sh_ddr_rready),
    .sh_cl_ddr_is_ready(sh_cl_ddr_is_ready),
    .cl_sh_apppf_irq_req(cl_sh_apppf_irq_req),
    .sh_cl_apppf_irq_ack(sh_cl_apppf_irq_ack),
    .sh_cl_dma_pcis_awid(sh_cl_dma_pcis_awid),
    .sh_cl_dma_pcis_awaddr(sh_cl_dma_pcis_awaddr),
    .sh_cl_dma_pcis_awlen(sh_cl_dma_pcis_awlen),
    .sh_cl_dma_pcis_awsize(sh_cl_dma_pcis_awsize),
    .sh_cl_dma_pcis_awvalid(sh_cl_dma_pcis_awvalid),
    .cl_sh_dma_pcis_awready(cl_sh_dma_pcis_awready),
    .sh_cl_dma_pcis_wdata(sh_cl_dma_pcis_wdata),
    .sh_cl_dma_pcis_wstrb(sh_cl_dma_pcis_wstrb),
    .sh_cl_dma_pcis_wlast(sh_cl_dma_pcis_wlast),
    .sh_cl_dma_pcis_wvalid(sh_cl_dma_pcis_wvalid),
    .cl_sh_dma_pcis_wready(cl_sh_dma_pcis_wready),
    .cl_sh_dma_pcis_bid(cl_sh_dma_pcis_bid),
    .cl_sh_dma_pcis_bresp(cl_sh_dma_pcis_bresp),
    .cl_sh_dma_pcis_bvalid(cl_sh_dma_pcis_bvalid),
    .sh_cl_dma_pcis_bready(sh_cl_dma_pcis_bready),
    .sh_cl_dma_pcis_arid(sh_cl_dma_pcis_arid),
    .sh_cl_dma_pcis_araddr(sh_cl_dma_pcis_araddr),
    .sh_cl_dma_pcis_arlen(sh_cl_dma_pcis_arlen),
    .sh_cl_dma_pcis_arsize(sh_cl_dma_pcis_arsize),
    .sh_cl_dma_pcis_arvalid(sh_cl_dma_pcis_arvalid),
    .cl_sh_dma_pcis_arready(cl_sh_dma_pcis_arready),
    .cl_sh_dma_pcis_rid(cl_sh_dma_pcis_rid),
    .cl_sh_dma_pcis_rdata(cl_sh_dma_pcis_rdata),
    .cl_sh_dma_pcis_rresp(cl_sh_dma_pcis_rresp),
    .cl_sh_dma_pcis_rlast(cl_sh_dma_pcis_rlast),
    .cl_sh_dma_pcis_rvalid(cl_sh_dma_pcis_rvalid),
    .sh_cl_dma_pcis_rready(sh_cl_dma_pcis_rready),
    .sda_cl_awvalid(sda_cl_awvalid),
    .sda_cl_awaddr(sda_cl_awaddr),
    .cl_sda_awready(cl_sda_awready),
    .sda_cl_wvalid(sda_cl_wvalid),
    .sda_cl_wdata(sda_cl_wdata),
    .sda_cl_wstrb(sda_cl_wstrb),
    .cl_sda_wready(cl_sda_wready),
    .cl_sda_bvalid(cl_sda_bvalid),
    .cl_sda_bresp(cl_sda_bresp),
    .sda_cl_bready(sda_cl_bready),
    .sda_cl_arvalid(sda_cl_arvalid),
    .sda_cl_araddr(sda_cl_araddr),
    .cl_sda_arready(cl_sda_arready),
    .cl_sda_rvalid(cl_sda_rvalid),
    .cl_sda_rdata(cl_sda_rdata),
    .cl_sda_rresp(cl_sda_rresp),
    .sda_cl_rready(sda_cl_rready),
    .sh_ocl_awvalid(sh_ocl_awvalid),
    .sh_ocl_awaddr(sh_ocl_awaddr),
    .ocl_sh_awready(ocl_sh_awready),
    .sh_ocl_wvalid(sh_ocl_wvalid),
    .sh_ocl_wdata(sh_ocl_wdata),
    .sh_ocl_wstrb(sh_ocl_wstrb),
    .ocl_sh_wready(ocl_sh_wready),
    .ocl_sh_bvalid(ocl_sh_bvalid),
    .ocl_sh_bresp(ocl_sh_bresp),
    .sh_ocl_bready(sh_ocl_bready),
    .sh_ocl_arvalid(sh_ocl_arvalid),
    .sh_ocl_araddr(sh_ocl_araddr),
    .ocl_sh_arready(ocl_sh_arready),
    .ocl_sh_rvalid(ocl_sh_rvalid),
    .ocl_sh_rdata(ocl_sh_rdata),
    .ocl_sh_rresp(ocl_sh_rresp),
    .sh_ocl_rready(sh_ocl_rready),
    .sh_bar1_awvalid(sh_bar1_awvalid),
    .sh_bar1_awaddr(sh_bar1_awaddr),
    .bar1_sh_awready(bar1_sh_awready),
    .sh_bar1_wvalid(sh_bar1_wvalid),
    .sh_bar1_wdata(sh_bar1_wdata),
    .sh_bar1_wstrb(sh_bar1_wstrb),
    .bar1_sh_wready(bar1_sh_wready),
    .bar1_sh_bvalid(bar1_sh_bvalid),
    .bar1_sh_bresp(bar1_sh_bresp),
    .sh_bar1_bready(sh_bar1_bready),
    .sh_bar1_arvalid(sh_bar1_arvalid),
    .sh_bar1_araddr(sh_bar1_araddr),
    .bar1_sh_arready(bar1_sh_arready),
    .bar1_sh_rvalid(bar1_sh_rvalid),
    .bar1_sh_rdata(bar1_sh_rdata),
    .bar1_sh_rresp(bar1_sh_rresp),
    .sh_bar1_rready(sh_bar1_rready),
    .drck(drck),
    .shift(shift),
    .update(update),
    .sel(sel),
    .runtest(runtest),
    .reset(reset),
    .capture(capture),
    .bscanid_en(bscanid_en),
    .sh_cl_glcount0(sh_cl_glcount0),
    .sh_cl_glcount1(sh_cl_glcount1)
	);
endmodule
