module IOBUF (
		output wire [0:0] dataout, //   dout.export
		input  wire [0:0] datain,  //    din.export
		input  wire [0:0] oe,      //     oe.export
		inout  wire [0:0] padio    // pad_io.export
	);
endmodule

